----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    16:44:11 03/21/2017 
-- Design Name: 
-- Module Name:    Adder - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.std_logic_unsigned.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Adder is
    Port ( OP1 : in  STD_LOGIC_Vector(31 downto 0);
           OP2 : in  STD_LOGIC_Vector(31 downto 0);
           RESULT : out  STD_LOGIC_Vector(31 downto 0));
end Adder;

architecture Behavioral of Adder is

	signal Result_aux : STD_LOGIC_VECTOR(31 downto 0) := (others => '0');

begin
	process(OP1,OP2)
	begin
		Result_aux <= OP1 + OP2;
	end process;
	
	RESULT <= Result_aux;
end Behavioral;

